// created by ivy on 2021/6/30

module Add (
    input [31:0] a,
    input [31:0] b,
    output [31:0] out
);
    // TO DO
    // use ~, !, |, & to implement an 32-bits adder
    // If the digits overflow, discard the overflow digits directly

endmodule
