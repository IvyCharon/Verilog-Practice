// created by ivy on 2021/6/30

module Add (
    input [31:0] a,
    input [31:0] b,
    output reg [31:0] sum
);
    // TO DO
    // use ^, !, ~, & to implement an 32-bits adder
    // If the digits overflow, discard the overflow digits directly

endmodule
