module zdo (
    input wire rst
);
    // TO DO
    
endmodule